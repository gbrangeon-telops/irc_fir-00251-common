----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 04/10/2024 11:25:32 AM
-- Design Name: 
-- Module Name: pgm_builder - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

library WORK;
use WORK.TEL2000.ALL;
use WORK.PROXY_DEFINE.ALL;

library STD;
use STD.TEXTIO.ALL;

entity pgm_builder is
    Generic (
        FILEPATH : string := "frame.pgm"
    );
    Port (
        clock  : in std_logic;
        data   : in t_axi4_stream_mosi128;
        config : in fpa_intf_cfg_type
    );
end pgm_builder;

architecture Behavioral of pgm_builder is
    file pgm : text;
begin

    process
    begin
        wait until rising_edge(clock) and data.tvalid = '1';
        
        file_open(pgm, FILEPATH, WRITE_MODE);
        
        write(pgm, "P2" & LF);
        write(pgm, "# Generated by pgm_builder" & LF);
        write(pgm, integer'image(to_integer(config.width)) & " " & integer'image(to_integer(config.height)) & LF);
        write(pgm, "65535" & LF);
        
        for y in 1 to to_integer(config.height) loop
            for x in 1 to to_integer(config.width) / 8 loop
                write(pgm, integer'image(to_integer(unsigned(data.tdata( 15 downto   0)))) & " ");
                write(pgm, integer'image(to_integer(unsigned(data.tdata( 31 downto  16)))) & " ");
                write(pgm, integer'image(to_integer(unsigned(data.tdata( 47 downto  32)))) & " ");
                write(pgm, integer'image(to_integer(unsigned(data.tdata( 63 downto  48)))) & " ");
                write(pgm, integer'image(to_integer(unsigned(data.tdata( 79 downto  64)))) & " ");
                write(pgm, integer'image(to_integer(unsigned(data.tdata( 95 downto  80)))) & " ");
                write(pgm, integer'image(to_integer(unsigned(data.tdata(111 downto  96)))) & " ");
                write(pgm, integer'image(to_integer(unsigned(data.tdata(127 downto 112)))) & " ");
                
                if data.tlast = '0' then
                    wait until rising_edge(clock) and data.tvalid = '1';
                end if;
            end loop;
            write(pgm, "" & LF);
        end loop;
        
        file_close(pgm);
    end process;

end Behavioral;
