-------------------------------------------------------------------------------
--
-- Title       : USART_TO_AXIS
-- Design      : Usart_tb
-- Author      : 
-- Company     : 
--
-------------------------------------------------------------------------------
--
-- File        : D:\Telops\FIR-00251-Common\VHDL\USART_B\sims\src\USART_TO_AXIS.vhd
-- Generated   : Fri Oct  9 11:49:23 2015
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {USART_TO_AXIS} architecture {USART_TO_AXIS}}

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity USART_TO_AXIS is
end USART_TO_AXIS;

--}} End of automatically maintained section

architecture USART_TO_AXIS of USART_TO_AXIS is
begin

	 -- enter your statements here --

end USART_TO_AXIS;
